Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.std_logic_unsigned.all;
Use IEEE.std_logic_arith.all;
Use work.mis_componentes.all;
---------------------------------------------------------------------------------------------------------
ENTITY MATRIZ_PARQUEADERO IS
PORT(	START: 				In std_logic;
		INGRESAR: 			In std_logic;
		SALIR: 				In std_logic;
		COD_AUTO_SALIDA: 	In std_logic_vector(3 downto 0);
		RESET: 				In std_logic;
		CLOCK: 				In std_logic;
		CLOCK_1Hz: 			In std_logic;
		CLOCK_100Hz:		In std_logic;
		
		DIRECCION_RAM:		Out std_logic_vector(3 downto 0);
		CONTENIDO_RAM:		Out std_logic;
		
		ENTRADA: 			Out std_logic;
		SALIDA: 				Out std_logic;
		DENEGADO: 			Out std_logic;
		COLUMNA_MATRIZ:	Out std_logic_vector(3 downto 0);
		FILA_MATRIZ:		Out std_logic_vector(3 downto 0);
		COLUMNA_LIB:		Out std_logic_vector(6 downto 0);
		FILA_LIB:			Out std_logic_vector(6 downto 0);
		DEC_P_LIBRES:		Out std_logic_vector(6 downto 0);
		UNID_P_LIBRES:		Out std_logic_vector(6 downto 0));
END MATRIZ_PARQUEADERO; 
---------------------------------------------------------------------------------------------------------
ARCHITECTURE estructural OF MATRIZ_PARQUEADERO IS
-------------------------------------------------------------------------------------------------------------
TYPE ESTADO IS (T0, T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16);
SIGNAL Y: ESTADO;

SIGNAL EN_CONT_DIRECC, RESET_CONT_DIRECC: std_logic;
SIGNAL DIRECCION: std_logic_vector(3 downto 0);
SIGNAL UNO_CERO: std_logic_vector(1 downto 0);
SIGNAL OCUPADO: std_logic;
SIGNAL WR: std_logic;
SIGNAL ADDRESS_RAM: std_logic_vector(3 downto 0);
SIGNAL CARRO_SALIDA: std_logic;
SIGNAL EN_TIME, RESET_TIME, IG_3SEG: std_logic;
SIGNAL TIME_PARPADEO: std_logic_vector(1 downto 0);
SIGNAL EN_CONT_LIBRES, LOAD_CONT_LIBRES, SUMA_PL, RESTA_PL, RESET_CONT_LIBRES, HAY_LIBRES: std_logic;
SIGNAL P_LIBRES: std_logic_vector(4 downto 0);
SIGNAL FF1, FF2, FF3, FF4, FF5, FF6, FF7, FF8, FF9, FF10, FF11, FF12, FF13, FF14, FF15, FF16: std_logic;
SIGNAL EN_FF, RESET_FF, RESET_M: std_logic;
SIGNAL P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16: std_logic;
SIGNAL TIME_FF, TIMEFF1, TIMEFF2, TIMEFF3, TIMEFF4, TIMEFF5, TIMEFF6, TIMEFF7, TIMEFF8, TIMEFF9, TIMEFF10, TIMEFF11, TIMEFF12, TIMEFF13, TIMEFF14, TIMEFF15, TIMEFF16: std_logic_vector(5 downto 0);
SIGNAL UN_MINUTO: std_logic;
SIGNAL COLUMN_0, COLUMN_1, COLUMN_2, COLUMN_3: std_logic_vector(3 downto 0);
SIGNAL EN_CONT_COLUMN, RESET_CONT_COLUMN: std_logic;
SIGNAL COLUMN_ACTIV: std_logic_vector(1 downto 0);
SIGNAL EN_MATRIZ, C0_ON, C1_ON, C2_ON, C3_ON: std_logic;
SIGNAL APAGAR_1, APAGAR_2: std_logic;
SIGNAL DEC_BCD_P_LIB, UNID_BCD_P_LIB: std_logic_vector(3 downto 0);
SIGNAL COLUMNA_BCD, FILA_BCD: std_logic_vector(3 downto 0);
SIGNAL SIN_USO_0, SIN_USO_1, SIN_USO_2: std_logic;
-------------------------------------------------------------------------------------------------------------
BEGIN
	MSS_TRANSICIONES: PROCESS(RESET, CLOCK)
	BEGIN
		IF RESET='1' THEN Y <= T0;
		ELSIF (CLOCK'EVENT AND CLOCK='1') THEN
			CASE Y IS
				WHEN T0 => IF START='0' THEN Y<=T0; ELSE Y<=T1; END IF;
				WHEN T1 => IF START='1' THEN Y<=T1; ELSE Y<=T2; END IF;
				WHEN T2 => IF (INGRESAR='0' AND SALIR='1') THEN Y<=T3;
							  ELSIF (INGRESAR='1' AND HAY_LIBRES='1') THEN Y<=T10;
							  ELSE Y<=T2; END IF;
				WHEN T3 => IF SALIR='0' THEN Y<=T4; ELSE Y<=T3; END IF;
				WHEN T4 => IF OCUPADO='0' THEN Y<=T2;
							  ELSIF UN_MINUTO='0' THEN Y<=T5;
							  ELSE Y<=T7; END IF;
				WHEN T5 => IF IG_3SEG='1' THEN Y<=T6; ELSE Y<=T5; END IF;
				WHEN T6 => Y<=T2;
				WHEN T7 => Y<=T8;
				WHEN T8 => IF IG_3SEG='1' THEN Y<=T6; ELSE Y<=T9; END IF;
				WHEN T9 => Y<=T8;
				WHEN T10 => IF INGRESAR='0' THEN Y<=T11; ELSE Y<=T10; END IF;
				WHEN T11 => IF OCUPADO='1' THEN Y<=T12; ELSE Y<=T13; END IF;
				WHEN T12 => Y<=T16;
				WHEN T13 => Y<=T14;
				WHEN T14 => IF IG_3SEG='1' THEN Y<=T6; ELSE Y<=T15; END IF;
				WHEN T15 => Y<=T14;
				WHEN T16 => Y<=T11;
			END CASE;
		END IF;
	END PROCESS;
	
	MSS_SALIDAS: PROCESS(Y, START, INGRESAR, SALIR, OCUPADO, IG_3SEG, HAY_LIBRES, UN_MINUTO)
	BEGIN
		APAGAR_1<='0'; APAGAR_2<='0'; ENTRADA<='0'; SALIDA<='0'; DENEGADO<='0'; 
		EN_CONT_DIRECC<='0'; RESET_CONT_DIRECC<='0'; 
		CARRO_SALIDA<='0'; UNO_CERO(0)<='0'; WR<='0'; 
		EN_TIME<='0'; RESET_TIME<='0'; 
		EN_CONT_LIBRES<='0'; RESET_CONT_LIBRES<='0'; LOAD_CONT_LIBRES<='0'; SUMA_PL<='0'; RESTA_PL<='0';
		EN_FF<='0'; RESET_FF<='0'; 
		EN_MATRIZ<='0'; RESET_M<='0'; EN_CONT_COLUMN<='0'; RESET_CONT_COLUMN<='0';
		
		
		CASE Y IS
			WHEN T0 =>  RESET_CONT_DIRECC<='1'; RESET_TIME<='1'; RESET_CONT_LIBRES<='1'; RESET_M<='1'; RESET_CONT_COLUMN<='1'; APAGAR_1<='1'; APAGAR_2<='1';
			WHEN T1 =>  RESET_CONT_DIRECC<='1'; RESET_TIME<='1'; RESET_M<='1'; RESET_CONT_COLUMN<='1'; APAGAR_1<='1'; APAGAR_2<='1';
							IF START='1' THEN RESET_CONT_LIBRES<='1'; ELSE EN_CONT_LIBRES<='1'; LOAD_CONT_LIBRES<='1'; END IF;
			WHEN T2 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1';
			WHEN T3 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1'; CARRO_SALIDA<='1';
			WHEN T4 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; CARRO_SALIDA<='1';
							IF OCUPADO='0' THEN APAGAR_2<='1'; END IF;
			WHEN T5 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; DENEGADO<='1'; EN_TIME<='1'; APAGAR_2<='1';
			WHEN T6 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; RESET_TIME<='1'; APAGAR_2<='1';
			WHEN T7 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; CARRO_SALIDA<='1'; WR<='1'; EN_CONT_LIBRES<='1'; SUMA_PL<='1'; RESET_FF<='1'; 
			WHEN T8 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; EN_TIME<='1'; SALIDA<='1'; CARRO_SALIDA<='1';
			WHEN T9 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; EN_TIME<='1'; CARRO_SALIDA<='1';
			WHEN T10 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1';
			WHEN T11 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1';
			WHEN T12 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1'; EN_CONT_DIRECC<='1';
			WHEN T13 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; UNO_CERO(0)<='1'; WR<='1'; EN_CONT_LIBRES<='1'; RESTA_PL<='1'; EN_FF<='1';
			WHEN T14 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; EN_TIME<='1'; ENTRADA<='1';
							 IF IG_3SEG='1' THEN RESET_CONT_DIRECC<='1'; APAGAR_2<='1'; END IF;
			WHEN T15 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; EN_TIME<='1';
			WHEN T16 =>  EN_MATRIZ<='1'; EN_CONT_COLUMN<='1'; APAGAR_2<='1';
		END CASE;
	END PROCESS;
	
	COLUMN_0 <= (NOT(P1) & NOT(P5) & NOT(P9) & NOT(P13));
	COLUMN_1 <= (NOT(P2) & NOT(P6) & NOT(P10) & NOT(P14));
	COLUMN_2 <= (NOT(P3) & NOT(P7) & NOT(P11) & NOT(P15));
	COLUMN_3 <= (NOT(P4) & NOT(P8) & NOT(P12) & NOT(P16));
	UNO_CERO(1) <= '0';
	FILA_MATRIZ <= (C0_ON & C1_ON & C2_ON & C3_ON);
	HAY_LIBRES <= (P_LIBRES(4) OR P_LIBRES(3) OR P_LIBRES(2) OR P_LIBRES(1) OR P_LIBRES(0));
	IG_3SEG <= (TIME_PARPADEO(1) AND TIME_PARPADEO(0));
	
	DIRECCION_RAM <= ADDRESS_RAM;
	CONTENIDO_RAM <= OCUPADO;
	
	CONTADOR_DIRECCIONES: CONTADOR_UP Port Map("0000", EN_CONT_DIRECC, '0', RESET_CONT_DIRECC, CLOCK, DIRECCION);
	--RAM_POSICIONES: RAM_PUESTOS Port Map(('0'&ADDRESS_RAM), CLOCK, UNO_CERO, WR, OCUPADO);
	MUX_RAM: MUX_16_1_bit Port Map(P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, ADDRESS_RAM, OCUPADO); 
	MUX1: MUX_2TO1 Port Map(DIRECCION, COD_AUTO_SALIDA, CARRO_SALIDA, ADDRESS_RAM); 
	CONTADOR_TIEMPO_PARPADEO: CONTADOR_UP_3bits Port Map("00", EN_TIME, '0', RESET_TIME, CLOCK_1Hz, TIME_PARPADEO);
	CONTADOR_POSICIONES_LIBRES: CONTADOR_UP_DOWN Port Map("10000", EN_CONT_LIBRES, LOAD_CONT_LIBRES, SUMA_PL, RESTA_PL, RESET_CONT_LIBRES, CLOCK, P_LIBRES);
	DEMULTIPLEXADOR: DEMUX_1TO16 Port Map('1', ADDRESS_RAM, FF1, FF2, FF3, FF4, FF5, FF6, FF7, FF8, FF9, FF10, FF11, FF12, FF13, FF14, FF15, FF16);
	PUESTO_1: FF_tipoD Port Map('1', (EN_FF AND FF1), ((FF1 AND RESET_FF) OR RESET_M), CLOCK, P1);
	CONTADOR_TIEMPO_P1: CONTADOR_UP_60LIM Port Map("000000", P1, '0', (NOT(P1)), CLOCK_1Hz, TIMEFF1); --1
	PUESTO_2: FF_tipoD Port Map('1', (EN_FF AND FF2), ((FF2 AND RESET_FF) OR RESET_M), CLOCK, P2);
	CONTADOR_TIEMPO_P2: CONTADOR_UP_60LIM Port Map("000000", P2, '0', (NOT(P2)), CLOCK_1Hz, TIMEFF2); --2
	PUESTO_3: FF_tipoD Port Map('1', (EN_FF AND FF3), ((FF3 AND RESET_FF) OR RESET_M), CLOCK, P3);
	CONTADOR_TIEMPO_P3: CONTADOR_UP_60LIM Port Map("000000", P3, '0', (NOT(P3)), CLOCK_1Hz, TIMEFF3); --3
	PUESTO_4: FF_tipoD Port Map('1', (EN_FF AND FF4), ((FF4 AND RESET_FF) OR RESET_M), CLOCK, P4);
	CONTADOR_TIEMPO_P4: CONTADOR_UP_60LIM Port Map("000000", P4, '0', (NOT(P4)), CLOCK_1Hz, TIMEFF4); --4
	PUESTO_5: FF_tipoD Port Map('1', (EN_FF AND FF5), ((FF5 AND RESET_FF) OR RESET_M), CLOCK, P5);
	CONTADOR_TIEMPO_P5: CONTADOR_UP_60LIM Port Map("000000", P5, '0', (NOT(P5)), CLOCK_1Hz, TIMEFF5); --5
	PUESTO_6: FF_tipoD Port Map('1', (EN_FF AND FF6), ((FF6 AND RESET_FF) OR RESET_M), CLOCK, P6);
	CONTADOR_TIEMPO_P6: CONTADOR_UP_60LIM Port Map("000000", P6, '0', (NOT(P6)), CLOCK_1Hz, TIMEFF6); --6
	PUESTO_7: FF_tipoD Port Map('1', (EN_FF AND FF7), ((FF7 AND RESET_FF) OR RESET_M), CLOCK, P7);
	CONTADOR_TIEMPO_P7: CONTADOR_UP_60LIM Port Map("000000", P7, '0', (NOT(P7)), CLOCK_1Hz, TIMEFF7); --7
	PUESTO_8: FF_tipoD Port Map('1', (EN_FF AND FF8), ((FF8 AND RESET_FF) OR RESET_M), CLOCK, P8);
	CONTADOR_TIEMPO_P8: CONTADOR_UP_60LIM Port Map("000000", P8, '0', (NOT(P8)), CLOCK_1Hz, TIMEFF8); --8
	PUESTO_9: FF_tipoD Port Map('1', (EN_FF AND FF9), ((FF9 AND RESET_FF) OR RESET_M), CLOCK, P9);
	CONTADOR_TIEMPO_P9: CONTADOR_UP_60LIM Port Map("000000", P9, '0', (NOT(P9)), CLOCK_1Hz, TIMEFF9); --9
	PUESTO_10: FF_tipoD Port Map('1', (EN_FF AND FF10), ((FF10 AND RESET_FF) OR RESET_M), CLOCK, P10);
	CONTADOR_TIEMPO_P10: CONTADOR_UP_60LIM Port Map("000000", P10, '0', (NOT(P10)), CLOCK_1Hz, TIMEFF10); --10
	PUESTO_11: FF_tipoD Port Map('1', (EN_FF AND FF11), ((FF11 AND RESET_FF) OR RESET_M), CLOCK, P11);
	CONTADOR_TIEMPO_P11: CONTADOR_UP_60LIM Port Map("000000", P11, '0', (NOT(P11)), CLOCK_1Hz, TIMEFF11); --11
	PUESTO_12: FF_tipoD Port Map('1', (EN_FF AND FF12), ((FF12 AND RESET_FF) OR RESET_M), CLOCK, P12);
	CONTADOR_TIEMPO_P12: CONTADOR_UP_60LIM Port Map("000000", P12, '0', (NOT(P12)), CLOCK_1Hz, TIMEFF12); --12
	PUESTO_13: FF_tipoD Port Map('1', (EN_FF AND FF13), ((FF13 AND RESET_FF) OR RESET_M), CLOCK, P13);
	CONTADOR_TIEMPO_P13: CONTADOR_UP_60LIM Port Map("000000", P13, '0', (NOT(P13)), CLOCK_1Hz, TIMEFF13); --13
	PUESTO_14: FF_tipoD Port Map('1', (EN_FF AND FF14), ((FF14 AND RESET_FF) OR RESET_M), CLOCK, P14);
	CONTADOR_TIEMPO_P14: CONTADOR_UP_60LIM Port Map("000000", P14, '0', (NOT(P14)), CLOCK_1Hz, TIMEFF14); --14
	PUESTO_15: FF_tipoD Port Map('1', (EN_FF AND FF15), ((FF15 AND RESET_FF) OR RESET_M), CLOCK, P15);
	CONTADOR_TIEMPO_P15: CONTADOR_UP_60LIM Port Map("000000", P15, '0', (NOT(P15)), CLOCK_1Hz, TIMEFF15); --15
	PUESTO_16: FF_tipoD Port Map('1', (EN_FF AND FF16), ((FF16 AND RESET_FF) OR RESET_M), CLOCK, P16);
	CONTADOR_TIEMPO_P16: CONTADOR_UP_60LIM Port Map("000000", P16, '0', (NOT(P16)), CLOCK_1Hz, TIMEFF16); --16
	MUX2: MUX_16_1 Port Map(TIMEFF1, TIMEFF2, TIMEFF3, TIMEFF4, TIMEFF5, TIMEFF6, TIMEFF7, TIMEFF8, TIMEFF9, TIMEFF10, TIMEFF11, TIMEFF12, TIMEFF13, TIMEFF14, TIMEFF15, TIMEFF16, ADDRESS_RAM, TIME_FF); 
	COMPARADOR_AL_MENOS_1_MIN: COMPARADOR Port Map(TIME_FF, "111100", SIN_USO_1, UN_MINUTO, SIN_USO_2);
	CONTADOR_ACTIVA_FILA: CONTADOR_UP_3bits Port Map("00", EN_CONT_COLUMN, '0', RESET_CONT_COLUMN, CLOCK_100Hz, COLUMN_ACTIV);
	COMPARADOR_FILA_ACTIVA: COMPARADOR_0to3 Port Map(COLUMN_ACTIV, EN_MATRIZ, C0_ON, C1_ON, C2_ON, C3_ON);
	MUX3: MUX_4_1 Port Map(COLUMN_0, COLUMN_1, COLUMN_2, COLUMN_3, EN_MATRIZ, COLUMN_ACTIV, COLUMNA_MATRIZ);
	BINARIO_A_BCD: DECODER_BINARIO_BCD Port Map(P_LIBRES, DEC_BCD_P_LIB, UNID_BCD_P_LIB);
	MUESTRA_POSICION_FORMATO_XY: POSICION_COLUM_FIL Port Map(ADDRESS_RAM, (NOT(APAGAR_2)), COLUMNA_BCD, FILA_BCD);
	DECENAS_PUESTOS_LIBRES: DECODER_7SEG Port Map(DEC_BCD_P_LIB, APAGAR_1, DEC_P_LIBRES);
	UNIDADES_PUESTOS_LIBRES: DECODER_7SEG Port Map(UNID_BCD_P_LIB, APAGAR_1, UNID_P_LIBRES);
	Y_COLUMNA: DECODER_7SEG Port Map(COLUMNA_BCD, APAGAR_2, COLUMNA_LIB);
	X_FILA: DECODER_7SEG Port Map(FILA_BCD, APAGAR_2, FILA_LIB);
	
END estructural;


	